.SUBCKT ActorSubckt NNIN1 NNIN2 NNIN3 NNIN4 NNIN5 NNIN6 NNIN7 NNIN8 NNIN9 NNIN10 NNIN11 NNIN12 NNIN13 NNIN14 NNIN15 NNIN16 NNIN17 NNIN18 NNIN19 NNOUT1

* LAYER 1: LINEAR
B1_1 L1_1 0 V=(V(NNIN1)*(-0.187835)+V(NNIN2)*(0.197037)+V(NNIN3)*(0.151082)+V(NNIN4)*(-0.188686)+V(NNIN5)*(-0.018063)+V(NNIN6)*(0.346796)+V(NNIN7)*(0.356271)+V(NNIN8)*(0.264235)+V(NNIN9)*(0.364792)+V(NNIN10)*(0.057384)+V(NNIN11)*(-0.215700)+V(NNIN12)*(-0.213923)+V(NNIN13)*(-0.011413)+V(NNIN14)*(0.209859)+V(NNIN15)*(0.129426)+V(NNIN16)*(-0.137232)+V(NNIN17)*(-0.133878)+V(NNIN18)*(-0.046964)+V(NNIN19)*(-0.089839)+(0.012259))
B1_2 L1_2 0 V=(V(NNIN1)*(-0.025406)+V(NNIN2)*(-0.059593)+V(NNIN3)*(0.074291)+V(NNIN4)*(0.148024)+V(NNIN5)*(-0.228714)+V(NNIN6)*(-0.370784)+V(NNIN7)*(-0.437327)+V(NNIN8)*(-0.499735)+V(NNIN9)*(-0.471179)+V(NNIN10)*(-0.353878)+V(NNIN11)*(-0.172490)+V(NNIN12)*(0.184754)+V(NNIN13)*(0.006535)+V(NNIN14)*(-0.160236)+V(NNIN15)*(0.022747)+V(NNIN16)*(-0.014039)+V(NNIN17)*(0.249059)+V(NNIN18)*(0.114698)+V(NNIN19)*(-0.033166)+(0.041824))
B1_3 L1_3 0 V=(V(NNIN1)*(-0.194591)+V(NNIN2)*(0.222355)+V(NNIN3)*(0.026852)+V(NNIN4)*(-0.070988)+V(NNIN5)*(-0.031901)+V(NNIN6)*(-0.081780)+V(NNIN7)*(0.218689)+V(NNIN8)*(-0.043062)+V(NNIN9)*(0.161831)+V(NNIN10)*(0.085902)+V(NNIN11)*(-0.026953)+V(NNIN12)*(0.078505)+V(NNIN13)*(0.032527)+V(NNIN14)*(-0.107019)+V(NNIN15)*(-0.035470)+V(NNIN16)*(0.198516)+V(NNIN17)*(0.039745)+V(NNIN18)*(0.141162)+V(NNIN19)*(0.098915)+(-0.060896))
B1_4 L1_4 0 V=(V(NNIN1)*(-0.032394)+V(NNIN2)*(-0.098517)+V(NNIN3)*(0.116745)+V(NNIN4)*(-0.025774)+V(NNIN5)*(0.028290)+V(NNIN6)*(-0.293050)+V(NNIN7)*(-0.573034)+V(NNIN8)*(-0.618205)+V(NNIN9)*(-0.550662)+V(NNIN10)*(-0.109252)+V(NNIN11)*(0.135085)+V(NNIN12)*(-0.060005)+V(NNIN13)*(0.126246)+V(NNIN14)*(-0.001368)+V(NNIN15)*(-0.217449)+V(NNIN16)*(0.266364)+V(NNIN17)*(-0.009185)+V(NNIN18)*(0.198671)+V(NNIN19)*(-0.064513)+(0.078688))
B1_5 L1_5 0 V=(V(NNIN1)*(-0.021998)+V(NNIN2)*(0.054118)+V(NNIN3)*(0.179899)+V(NNIN4)*(0.013463)+V(NNIN5)*(0.208443)+V(NNIN6)*(0.338851)+V(NNIN7)*(0.247920)+V(NNIN8)*(0.060406)+V(NNIN9)*(0.224639)+V(NNIN10)*(0.060214)+V(NNIN11)*(-0.012066)+V(NNIN12)*(-0.181457)+V(NNIN13)*(0.110913)+V(NNIN14)*(0.006647)+V(NNIN15)*(0.051852)+V(NNIN16)*(0.111980)+V(NNIN17)*(0.024182)+V(NNIN18)*(0.108002)+V(NNIN19)*(0.108678)+(-0.055250))
B1_6 L1_6 0 V=(V(NNIN1)*(0.243712)+V(NNIN2)*(-0.023402)+V(NNIN3)*(0.061606)+V(NNIN4)*(0.121012)+V(NNIN5)*(0.071321)+V(NNIN6)*(-0.440299)+V(NNIN7)*(-0.350028)+V(NNIN8)*(-0.213697)+V(NNIN9)*(-0.257951)+V(NNIN10)*(-0.402929)+V(NNIN11)*(0.170346)+V(NNIN12)*(0.048290)+V(NNIN13)*(-0.187791)+V(NNIN14)*(0.164198)+V(NNIN15)*(-0.177652)+V(NNIN16)*(0.049732)+V(NNIN17)*(0.043303)+V(NNIN18)*(0.027413)+V(NNIN19)*(-0.214475)+(0.143684))
B1_7 L1_7 0 V=(V(NNIN1)*(0.051206)+V(NNIN2)*(0.167387)+V(NNIN3)*(-0.045525)+V(NNIN4)*(-0.156498)+V(NNIN5)*(-0.228754)+V(NNIN6)*(0.111369)+V(NNIN7)*(0.011999)+V(NNIN8)*(0.200927)+V(NNIN9)*(0.151962)+V(NNIN10)*(-0.166789)+V(NNIN11)*(0.219529)+V(NNIN12)*(0.190513)+V(NNIN13)*(-0.104399)+V(NNIN14)*(-0.174903)+V(NNIN15)*(-0.004463)+V(NNIN16)*(-0.185371)+V(NNIN17)*(0.094402)+V(NNIN18)*(0.008410)+V(NNIN19)*(0.094985)+(-0.150895))
B1_8 L1_8 0 V=(V(NNIN1)*(0.132044)+V(NNIN2)*(0.042355)+V(NNIN3)*(-0.000638)+V(NNIN4)*(-0.137456)+V(NNIN5)*(0.071250)+V(NNIN6)*(-0.326733)+V(NNIN7)*(-0.623109)+V(NNIN8)*(-0.522577)+V(NNIN9)*(-0.359460)+V(NNIN10)*(-0.329283)+V(NNIN11)*(0.208018)+V(NNIN12)*(0.223389)+V(NNIN13)*(0.189608)+V(NNIN14)*(-0.132802)+V(NNIN15)*(-0.224808)+V(NNIN16)*(0.068102)+V(NNIN17)*(-0.137348)+V(NNIN18)*(0.336230)+V(NNIN19)*(-0.224338)+(-0.113574))
B1_9 L1_9 0 V=(V(NNIN1)*(0.145281)+V(NNIN2)*(-0.147393)+V(NNIN3)*(-0.092598)+V(NNIN4)*(0.104402)+V(NNIN5)*(-0.171596)+V(NNIN6)*(-0.139623)+V(NNIN7)*(-0.412102)+V(NNIN8)*(0.023180)+V(NNIN9)*(-0.182356)+V(NNIN10)*(-0.229485)+V(NNIN11)*(-0.103287)+V(NNIN12)*(0.007527)+V(NNIN13)*(-0.006712)+V(NNIN14)*(0.108541)+V(NNIN15)*(-0.139685)+V(NNIN16)*(0.046694)+V(NNIN17)*(-0.003202)+V(NNIN18)*(0.025280)+V(NNIN19)*(0.002795)+(0.179033))
B1_10 L1_10 0 V=(V(NNIN1)*(0.070409)+V(NNIN2)*(0.164033)+V(NNIN3)*(0.244572)+V(NNIN4)*(-0.029037)+V(NNIN5)*(0.188169)+V(NNIN6)*(-0.345411)+V(NNIN7)*(-0.590108)+V(NNIN8)*(-0.401725)+V(NNIN9)*(-0.384498)+V(NNIN10)*(-0.130841)+V(NNIN11)*(0.053141)+V(NNIN12)*(0.102015)+V(NNIN13)*(0.210297)+V(NNIN14)*(0.192123)+V(NNIN15)*(0.168676)+V(NNIN16)*(0.174673)+V(NNIN17)*(0.247487)+V(NNIN18)*(0.073448)+V(NNIN19)*(-0.043875)+(0.009236))
B1_11 L1_11 0 V=(V(NNIN1)*(0.018580)+V(NNIN2)*(0.106152)+V(NNIN3)*(-0.146703)+V(NNIN4)*(-0.050215)+V(NNIN5)*(0.151428)+V(NNIN6)*(-0.027647)+V(NNIN7)*(-0.071436)+V(NNIN8)*(-0.039814)+V(NNIN9)*(-0.117572)+V(NNIN10)*(0.154143)+V(NNIN11)*(-0.220481)+V(NNIN12)*(-0.218456)+V(NNIN13)*(0.178891)+V(NNIN14)*(-0.167114)+V(NNIN15)*(-0.055060)+V(NNIN16)*(0.157647)+V(NNIN17)*(0.046717)+V(NNIN18)*(0.103013)+V(NNIN19)*(0.149165)+(0.010630))
B1_12 L1_12 0 V=(V(NNIN1)*(0.111196)+V(NNIN2)*(0.163189)+V(NNIN3)*(0.017679)+V(NNIN4)*(-0.120619)+V(NNIN5)*(0.139055)+V(NNIN6)*(-0.477833)+V(NNIN7)*(-0.319011)+V(NNIN8)*(-0.483203)+V(NNIN9)*(-0.137387)+V(NNIN10)*(-0.024143)+V(NNIN11)*(0.058294)+V(NNIN12)*(0.078836)+V(NNIN13)*(-0.113483)+V(NNIN14)*(0.065485)+V(NNIN15)*(-0.212244)+V(NNIN16)*(0.195776)+V(NNIN17)*(0.110271)+V(NNIN18)*(0.160766)+V(NNIN19)*(-0.236357)+(0.139979))
B1_13 L1_13 0 V=(V(NNIN1)*(0.197333)+V(NNIN2)*(0.071427)+V(NNIN3)*(-0.159528)+V(NNIN4)*(0.050005)+V(NNIN5)*(0.098089)+V(NNIN6)*(-0.264113)+V(NNIN7)*(-0.221473)+V(NNIN8)*(-0.257759)+V(NNIN9)*(-0.062113)+V(NNIN10)*(-0.331873)+V(NNIN11)*(0.185680)+V(NNIN12)*(0.017311)+V(NNIN13)*(0.093073)+V(NNIN14)*(-0.264433)+V(NNIN15)*(-0.013742)+V(NNIN16)*(-0.022265)+V(NNIN17)*(0.121856)+V(NNIN18)*(0.247234)+V(NNIN19)*(-0.212221)+(-0.181094))
B1_14 L1_14 0 V=(V(NNIN1)*(0.092795)+V(NNIN2)*(-0.131451)+V(NNIN3)*(0.067784)+V(NNIN4)*(0.199867)+V(NNIN5)*(0.083467)+V(NNIN6)*(-0.085962)+V(NNIN7)*(0.006086)+V(NNIN8)*(0.137580)+V(NNIN9)*(0.091494)+V(NNIN10)*(-0.201919)+V(NNIN11)*(0.005372)+V(NNIN12)*(0.119953)+V(NNIN13)*(-0.240166)+V(NNIN14)*(0.137284)+V(NNIN15)*(-0.075683)+V(NNIN16)*(-0.042859)+V(NNIN17)*(-0.022134)+V(NNIN18)*(0.215906)+V(NNIN19)*(0.185883)+(0.057750))
B1_15 L1_15 0 V=(V(NNIN1)*(0.185694)+V(NNIN2)*(0.160021)+V(NNIN3)*(-0.174112)+V(NNIN4)*(-0.026573)+V(NNIN5)*(-0.029825)+V(NNIN6)*(0.082142)+V(NNIN7)*(-0.113534)+V(NNIN8)*(0.190097)+V(NNIN9)*(0.057834)+V(NNIN10)*(0.089089)+V(NNIN11)*(-0.162961)+V(NNIN12)*(0.079286)+V(NNIN13)*(-0.138237)+V(NNIN14)*(-0.079237)+V(NNIN15)*(-0.154167)+V(NNIN16)*(-0.119913)+V(NNIN17)*(0.226834)+V(NNIN18)*(-0.113172)+V(NNIN19)*(0.244854)+(-0.095164))
B1_16 L1_16 0 V=(V(NNIN1)*(-0.239539)+V(NNIN2)*(-0.098096)+V(NNIN3)*(0.190766)+V(NNIN4)*(-0.082242)+V(NNIN5)*(-0.198098)+V(NNIN6)*(0.131174)+V(NNIN7)*(-0.161442)+V(NNIN8)*(0.007068)+V(NNIN9)*(0.058327)+V(NNIN10)*(0.149326)+V(NNIN11)*(0.023621)+V(NNIN12)*(-0.090088)+V(NNIN13)*(-0.011613)+V(NNIN14)*(-0.155141)+V(NNIN15)*(0.124846)+V(NNIN16)*(-0.209904)+V(NNIN17)*(0.039911)+V(NNIN18)*(0.082288)+V(NNIN19)*(0.039236)+(0.184598))
B1_17 L1_17 0 V=(V(NNIN1)*(0.120431)+V(NNIN2)*(0.022086)+V(NNIN3)*(-0.124898)+V(NNIN4)*(0.130928)+V(NNIN5)*(-0.237651)+V(NNIN6)*(0.094930)+V(NNIN7)*(0.101692)+V(NNIN8)*(-0.247038)+V(NNIN9)*(0.122595)+V(NNIN10)*(-0.109562)+V(NNIN11)*(-0.114721)+V(NNIN12)*(0.015255)+V(NNIN13)*(-0.263123)+V(NNIN14)*(0.013987)+V(NNIN15)*(-0.122284)+V(NNIN16)*(0.154749)+V(NNIN17)*(-0.192076)+V(NNIN18)*(0.032642)+V(NNIN19)*(0.203884)+(-0.097527))
B1_18 L1_18 0 V=(V(NNIN1)*(-0.174099)+V(NNIN2)*(0.068771)+V(NNIN3)*(0.125779)+V(NNIN4)*(0.124408)+V(NNIN5)*(0.091522)+V(NNIN6)*(-0.357070)+V(NNIN7)*(-0.500270)+V(NNIN8)*(-0.184505)+V(NNIN9)*(-0.179154)+V(NNIN10)*(-0.051121)+V(NNIN11)*(0.301489)+V(NNIN12)*(0.075938)+V(NNIN13)*(-0.082657)+V(NNIN14)*(0.084193)+V(NNIN15)*(-0.220308)+V(NNIN16)*(0.108667)+V(NNIN17)*(-0.133203)+V(NNIN18)*(0.418510)+V(NNIN19)*(-0.107220)+(-0.172327))
B1_19 L1_19 0 V=(V(NNIN1)*(-0.166474)+V(NNIN2)*(-0.094571)+V(NNIN3)*(-0.202327)+V(NNIN4)*(0.141873)+V(NNIN5)*(0.128971)+V(NNIN6)*(-0.417669)+V(NNIN7)*(-0.456960)+V(NNIN8)*(-0.319429)+V(NNIN9)*(-0.496575)+V(NNIN10)*(-0.193563)+V(NNIN11)*(0.211374)+V(NNIN12)*(0.074342)+V(NNIN13)*(-0.068136)+V(NNIN14)*(-0.201151)+V(NNIN15)*(-0.174232)+V(NNIN16)*(0.232727)+V(NNIN17)*(0.050694)+V(NNIN18)*(0.026415)+V(NNIN19)*(-0.001912)+(0.300904))
B1_20 L1_20 0 V=(V(NNIN1)*(0.041959)+V(NNIN2)*(-0.221451)+V(NNIN3)*(0.035539)+V(NNIN4)*(0.096598)+V(NNIN5)*(0.143659)+V(NNIN6)*(0.557533)+V(NNIN7)*(0.504040)+V(NNIN8)*(0.533843)+V(NNIN9)*(0.398986)+V(NNIN10)*(0.091974)+V(NNIN11)*(-0.102297)+V(NNIN12)*(-0.157181)+V(NNIN13)*(0.112657)+V(NNIN14)*(-0.014067)+V(NNIN15)*(-0.157223)+V(NNIN16)*(-0.025557)+V(NNIN17)*(0.181386)+V(NNIN18)*(-0.327235)+V(NNIN19)*(-0.179674)+(-0.128325))
B1_21 L1_21 0 V=(V(NNIN1)*(-0.073658)+V(NNIN2)*(0.044392)+V(NNIN3)*(-0.046036)+V(NNIN4)*(0.154099)+V(NNIN5)*(0.213831)+V(NNIN6)*(-0.027227)+V(NNIN7)*(0.138493)+V(NNIN8)*(-0.100307)+V(NNIN9)*(-0.040434)+V(NNIN10)*(-0.245570)+V(NNIN11)*(0.224094)+V(NNIN12)*(-0.225704)+V(NNIN13)*(0.136245)+V(NNIN14)*(0.166757)+V(NNIN15)*(0.153984)+V(NNIN16)*(0.096344)+V(NNIN17)*(-0.210948)+V(NNIN18)*(0.026739)+V(NNIN19)*(0.199261)+(0.013101))
B1_22 L1_22 0 V=(V(NNIN1)*(0.216841)+V(NNIN2)*(0.157171)+V(NNIN3)*(-0.190266)+V(NNIN4)*(-0.205267)+V(NNIN5)*(-0.126539)+V(NNIN6)*(0.551522)+V(NNIN7)*(0.310737)+V(NNIN8)*(0.118020)+V(NNIN9)*(0.317833)+V(NNIN10)*(0.223076)+V(NNIN11)*(0.102043)+V(NNIN12)*(-0.050090)+V(NNIN13)*(-0.050611)+V(NNIN14)*(0.153168)+V(NNIN15)*(-0.058723)+V(NNIN16)*(-0.085094)+V(NNIN17)*(0.121964)+V(NNIN18)*(-0.407449)+V(NNIN19)*(-0.188163)+(0.015877))
B1_23 L1_23 0 V=(V(NNIN1)*(-0.024562)+V(NNIN2)*(-0.029706)+V(NNIN3)*(-0.050060)+V(NNIN4)*(0.129204)+V(NNIN5)*(0.047362)+V(NNIN6)*(0.395962)+V(NNIN7)*(0.578066)+V(NNIN8)*(0.212871)+V(NNIN9)*(0.355679)+V(NNIN10)*(0.307328)+V(NNIN11)*(-0.303775)+V(NNIN12)*(0.073000)+V(NNIN13)*(-0.134230)+V(NNIN14)*(-0.016408)+V(NNIN15)*(0.096736)+V(NNIN16)*(-0.209855)+V(NNIN17)*(-0.173504)+V(NNIN18)*(-0.177329)+V(NNIN19)*(-0.128202)+(0.009020))
B1_24 L1_24 0 V=(V(NNIN1)*(-0.124833)+V(NNIN2)*(0.040730)+V(NNIN3)*(0.280866)+V(NNIN4)*(0.297640)+V(NNIN5)*(-0.053797)+V(NNIN6)*(-0.281579)+V(NNIN7)*(-0.565173)+V(NNIN8)*(-0.567019)+V(NNIN9)*(-0.470249)+V(NNIN10)*(-0.368079)+V(NNIN11)*(0.165676)+V(NNIN12)*(0.133803)+V(NNIN13)*(-0.057974)+V(NNIN14)*(0.150044)+V(NNIN15)*(-0.046589)+V(NNIN16)*(-0.015215)+V(NNIN17)*(-0.068992)+V(NNIN18)*(0.185433)+V(NNIN19)*(-0.133465)+(-0.055445))
B1_25 L1_25 0 V=(V(NNIN1)*(-0.189934)+V(NNIN2)*(-0.071487)+V(NNIN3)*(-0.064349)+V(NNIN4)*(-0.241487)+V(NNIN5)*(0.065749)+V(NNIN6)*(0.617938)+V(NNIN7)*(0.430792)+V(NNIN8)*(0.440432)+V(NNIN9)*(0.247722)+V(NNIN10)*(0.175817)+V(NNIN11)*(-0.032976)+V(NNIN12)*(-0.235204)+V(NNIN13)*(0.221710)+V(NNIN14)*(0.226070)+V(NNIN15)*(0.061159)+V(NNIN16)*(0.183101)+V(NNIN17)*(-0.013486)+V(NNIN18)*(-0.055414)+V(NNIN19)*(-0.061706)+(-0.037907))
B1_26 L1_26 0 V=(V(NNIN1)*(0.055211)+V(NNIN2)*(0.174869)+V(NNIN3)*(0.074748)+V(NNIN4)*(-0.025610)+V(NNIN5)*(0.059403)+V(NNIN6)*(0.170629)+V(NNIN7)*(0.105821)+V(NNIN8)*(0.073712)+V(NNIN9)*(0.012435)+V(NNIN10)*(0.118489)+V(NNIN11)*(-0.111561)+V(NNIN12)*(0.195907)+V(NNIN13)*(0.062281)+V(NNIN14)*(0.055234)+V(NNIN15)*(-0.094286)+V(NNIN16)*(-0.023397)+V(NNIN17)*(-0.184330)+V(NNIN18)*(-0.033463)+V(NNIN19)*(0.206561)+(0.224040))
B1_27 L1_27 0 V=(V(NNIN1)*(0.200129)+V(NNIN2)*(0.135256)+V(NNIN3)*(-0.011541)+V(NNIN4)*(-0.215175)+V(NNIN5)*(-0.071305)+V(NNIN6)*(0.294306)+V(NNIN7)*(-0.081898)+V(NNIN8)*(0.005150)+V(NNIN9)*(-0.029904)+V(NNIN10)*(-0.087558)+V(NNIN11)*(-0.126490)+V(NNIN12)*(0.061601)+V(NNIN13)*(-0.161145)+V(NNIN14)*(0.209347)+V(NNIN15)*(0.004731)+V(NNIN16)*(0.074711)+V(NNIN17)*(0.170995)+V(NNIN18)*(-0.035691)+V(NNIN19)*(0.181768)+(0.078712))
B1_28 L1_28 0 V=(V(NNIN1)*(-0.029492)+V(NNIN2)*(0.208049)+V(NNIN3)*(-0.071291)+V(NNIN4)*(0.247687)+V(NNIN5)*(0.141239)+V(NNIN6)*(0.832952)+V(NNIN7)*(0.777020)+V(NNIN8)*(0.741771)+V(NNIN9)*(0.555968)+V(NNIN10)*(0.271659)+V(NNIN11)*(-0.189062)+V(NNIN12)*(-0.013367)+V(NNIN13)*(0.203361)+V(NNIN14)*(0.114993)+V(NNIN15)*(0.024905)+V(NNIN16)*(-0.086650)+V(NNIN17)*(0.062793)+V(NNIN18)*(-0.061211)+V(NNIN19)*(-0.072456)+(-0.181916))
B1_29 L1_29 0 V=(V(NNIN1)*(0.090402)+V(NNIN2)*(0.239014)+V(NNIN3)*(-0.014709)+V(NNIN4)*(0.131365)+V(NNIN5)*(-0.157683)+V(NNIN6)*(-0.320992)+V(NNIN7)*(-0.620720)+V(NNIN8)*(-0.516724)+V(NNIN9)*(-0.405574)+V(NNIN10)*(-0.431949)+V(NNIN11)*(0.102963)+V(NNIN12)*(-0.030251)+V(NNIN13)*(0.050984)+V(NNIN14)*(0.130764)+V(NNIN15)*(0.176403)+V(NNIN16)*(0.029301)+V(NNIN17)*(0.230754)+V(NNIN18)*(0.147824)+V(NNIN19)*(-0.205482)+(-0.036427))
B1_30 L1_30 0 V=(V(NNIN1)*(0.217882)+V(NNIN2)*(-0.085144)+V(NNIN3)*(0.226931)+V(NNIN4)*(-0.132610)+V(NNIN5)*(-0.195499)+V(NNIN6)*(0.098202)+V(NNIN7)*(-0.019104)+V(NNIN8)*(-0.179339)+V(NNIN9)*(-0.107424)+V(NNIN10)*(-0.135671)+V(NNIN11)*(-0.192866)+V(NNIN12)*(0.226814)+V(NNIN13)*(-0.037411)+V(NNIN14)*(0.100690)+V(NNIN15)*(0.056922)+V(NNIN16)*(-0.149713)+V(NNIN17)*(0.157482)+V(NNIN18)*(-0.195264)+V(NNIN19)*(0.153632)+(0.030606))
B1_31 L1_31 0 V=(V(NNIN1)*(0.102189)+V(NNIN2)*(-0.151753)+V(NNIN3)*(0.103470)+V(NNIN4)*(0.259002)+V(NNIN5)*(-0.127119)+V(NNIN6)*(-0.429983)+V(NNIN7)*(-0.504416)+V(NNIN8)*(-0.415815)+V(NNIN9)*(-0.550370)+V(NNIN10)*(-0.104822)+V(NNIN11)*(0.042265)+V(NNIN12)*(0.093003)+V(NNIN13)*(-0.091625)+V(NNIN14)*(0.134023)+V(NNIN15)*(0.186064)+V(NNIN16)*(-0.082767)+V(NNIN17)*(0.207266)+V(NNIN18)*(0.045173)+V(NNIN19)*(-0.123871)+(0.042563))
B1_32 L1_32 0 V=(V(NNIN1)*(0.017329)+V(NNIN2)*(0.122072)+V(NNIN3)*(0.084277)+V(NNIN4)*(-0.069829)+V(NNIN5)*(0.004634)+V(NNIN6)*(0.280411)+V(NNIN7)*(-0.029350)+V(NNIN8)*(-0.050863)+V(NNIN9)*(0.245121)+V(NNIN10)*(0.219867)+V(NNIN11)*(0.126124)+V(NNIN12)*(-0.116348)+V(NNIN13)*(-0.137829)+V(NNIN14)*(-0.172825)+V(NNIN15)*(0.097314)+V(NNIN16)*(-0.044721)+V(NNIN17)*(0.148850)+V(NNIN18)*(-0.174395)+V(NNIN19)*(0.203672)+(0.099017))
* ACTIVATION LAYER 1: RELU
B_ACT1_1 L_ACT1_1 0 V=(IF(V(L1_1)>0,V(L1_1),0))
B_ACT1_2 L_ACT1_2 0 V=(IF(V(L1_2)>0,V(L1_2),0))
B_ACT1_3 L_ACT1_3 0 V=(IF(V(L1_3)>0,V(L1_3),0))
B_ACT1_4 L_ACT1_4 0 V=(IF(V(L1_4)>0,V(L1_4),0))
B_ACT1_5 L_ACT1_5 0 V=(IF(V(L1_5)>0,V(L1_5),0))
B_ACT1_6 L_ACT1_6 0 V=(IF(V(L1_6)>0,V(L1_6),0))
B_ACT1_7 L_ACT1_7 0 V=(IF(V(L1_7)>0,V(L1_7),0))
B_ACT1_8 L_ACT1_8 0 V=(IF(V(L1_8)>0,V(L1_8),0))
B_ACT1_9 L_ACT1_9 0 V=(IF(V(L1_9)>0,V(L1_9),0))
B_ACT1_10 L_ACT1_10 0 V=(IF(V(L1_10)>0,V(L1_10),0))
B_ACT1_11 L_ACT1_11 0 V=(IF(V(L1_11)>0,V(L1_11),0))
B_ACT1_12 L_ACT1_12 0 V=(IF(V(L1_12)>0,V(L1_12),0))
B_ACT1_13 L_ACT1_13 0 V=(IF(V(L1_13)>0,V(L1_13),0))
B_ACT1_14 L_ACT1_14 0 V=(IF(V(L1_14)>0,V(L1_14),0))
B_ACT1_15 L_ACT1_15 0 V=(IF(V(L1_15)>0,V(L1_15),0))
B_ACT1_16 L_ACT1_16 0 V=(IF(V(L1_16)>0,V(L1_16),0))
B_ACT1_17 L_ACT1_17 0 V=(IF(V(L1_17)>0,V(L1_17),0))
B_ACT1_18 L_ACT1_18 0 V=(IF(V(L1_18)>0,V(L1_18),0))
B_ACT1_19 L_ACT1_19 0 V=(IF(V(L1_19)>0,V(L1_19),0))
B_ACT1_20 L_ACT1_20 0 V=(IF(V(L1_20)>0,V(L1_20),0))
B_ACT1_21 L_ACT1_21 0 V=(IF(V(L1_21)>0,V(L1_21),0))
B_ACT1_22 L_ACT1_22 0 V=(IF(V(L1_22)>0,V(L1_22),0))
B_ACT1_23 L_ACT1_23 0 V=(IF(V(L1_23)>0,V(L1_23),0))
B_ACT1_24 L_ACT1_24 0 V=(IF(V(L1_24)>0,V(L1_24),0))
B_ACT1_25 L_ACT1_25 0 V=(IF(V(L1_25)>0,V(L1_25),0))
B_ACT1_26 L_ACT1_26 0 V=(IF(V(L1_26)>0,V(L1_26),0))
B_ACT1_27 L_ACT1_27 0 V=(IF(V(L1_27)>0,V(L1_27),0))
B_ACT1_28 L_ACT1_28 0 V=(IF(V(L1_28)>0,V(L1_28),0))
B_ACT1_29 L_ACT1_29 0 V=(IF(V(L1_29)>0,V(L1_29),0))
B_ACT1_30 L_ACT1_30 0 V=(IF(V(L1_30)>0,V(L1_30),0))
B_ACT1_31 L_ACT1_31 0 V=(IF(V(L1_31)>0,V(L1_31),0))
B_ACT1_32 L_ACT1_32 0 V=(IF(V(L1_32)>0,V(L1_32),0))
* LAYER 2: LINEAR
B2_1 L2_1 0 V=(V(L_ACT1_1)*(0.041032)+V(L_ACT1_2)*(-0.069925)+V(L_ACT1_3)*(-0.076361)+V(L_ACT1_4)*(0.168700)+V(L_ACT1_5)*(0.065466)+V(L_ACT1_6)*(0.032381)+V(L_ACT1_7)*(-0.010142)+V(L_ACT1_8)*(0.135234)+V(L_ACT1_9)*(0.092256)+V(L_ACT1_10)*(0.006393)+V(L_ACT1_11)*(0.014046)+V(L_ACT1_12)*(0.000266)+V(L_ACT1_13)*(-0.058433)+V(L_ACT1_14)*(0.132049)+V(L_ACT1_15)*(-0.158908)+V(L_ACT1_16)*(-0.072086)+V(L_ACT1_17)*(-0.073096)+V(L_ACT1_18)*(0.075029)+V(L_ACT1_19)*(0.109545)+V(L_ACT1_20)*(0.052473)+V(L_ACT1_21)*(0.067381)+V(L_ACT1_22)*(0.111823)+V(L_ACT1_23)*(0.085856)+V(L_ACT1_24)*(0.059757)+V(L_ACT1_25)*(0.007457)+V(L_ACT1_26)*(0.175136)+V(L_ACT1_27)*(-0.113008)+V(L_ACT1_28)*(-0.088805)+V(L_ACT1_29)*(0.053813)+V(L_ACT1_30)*(-0.134330)+V(L_ACT1_31)*(0.014576)+V(L_ACT1_32)*(-0.136416)+(-0.123922))
B2_2 L2_2 0 V=(V(L_ACT1_1)*(0.057110)+V(L_ACT1_2)*(-0.236621)+V(L_ACT1_3)*(0.105213)+V(L_ACT1_4)*(0.114241)+V(L_ACT1_5)*(0.085778)+V(L_ACT1_6)*(0.026632)+V(L_ACT1_7)*(-0.005471)+V(L_ACT1_8)*(-0.029184)+V(L_ACT1_9)*(-0.182234)+V(L_ACT1_10)*(-0.067689)+V(L_ACT1_11)*(0.028206)+V(L_ACT1_12)*(-0.150909)+V(L_ACT1_13)*(-0.135439)+V(L_ACT1_14)*(-0.094205)+V(L_ACT1_15)*(0.177017)+V(L_ACT1_16)*(0.055103)+V(L_ACT1_17)*(-0.085057)+V(L_ACT1_18)*(-0.083625)+V(L_ACT1_19)*(-0.156551)+V(L_ACT1_20)*(0.204790)+V(L_ACT1_21)*(0.152160)+V(L_ACT1_22)*(0.141543)+V(L_ACT1_23)*(0.129641)+V(L_ACT1_24)*(0.007440)+V(L_ACT1_25)*(0.086106)+V(L_ACT1_26)*(0.139288)+V(L_ACT1_27)*(-0.015487)+V(L_ACT1_28)*(0.354572)+V(L_ACT1_29)*(0.011251)+V(L_ACT1_30)*(-0.033577)+V(L_ACT1_31)*(0.148711)+V(L_ACT1_32)*(0.129275)+(0.127831))
B2_3 L2_3 0 V=(V(L_ACT1_1)*(-0.031306)+V(L_ACT1_2)*(-0.097893)+V(L_ACT1_3)*(0.118884)+V(L_ACT1_4)*(-0.062958)+V(L_ACT1_5)*(0.109945)+V(L_ACT1_6)*(-0.081889)+V(L_ACT1_7)*(0.085534)+V(L_ACT1_8)*(0.054618)+V(L_ACT1_9)*(-0.109858)+V(L_ACT1_10)*(0.076662)+V(L_ACT1_11)*(-0.088389)+V(L_ACT1_12)*(0.101939)+V(L_ACT1_13)*(-0.020884)+V(L_ACT1_14)*(-0.052981)+V(L_ACT1_15)*(0.113844)+V(L_ACT1_16)*(-0.003712)+V(L_ACT1_17)*(0.176262)+V(L_ACT1_18)*(-0.021857)+V(L_ACT1_19)*(-0.051013)+V(L_ACT1_20)*(0.185074)+V(L_ACT1_21)*(-0.037068)+V(L_ACT1_22)*(0.001533)+V(L_ACT1_23)*(0.191360)+V(L_ACT1_24)*(0.119628)+V(L_ACT1_25)*(0.026189)+V(L_ACT1_26)*(-0.052112)+V(L_ACT1_27)*(0.167044)+V(L_ACT1_28)*(0.100656)+V(L_ACT1_29)*(-0.118773)+V(L_ACT1_30)*(0.165408)+V(L_ACT1_31)*(0.031616)+V(L_ACT1_32)*(0.043423)+(-0.014603))
B2_4 L2_4 0 V=(V(L_ACT1_1)*(-0.210671)+V(L_ACT1_2)*(0.240926)+V(L_ACT1_3)*(-0.130949)+V(L_ACT1_4)*(0.019924)+V(L_ACT1_5)*(0.016914)+V(L_ACT1_6)*(-0.004464)+V(L_ACT1_7)*(-0.147269)+V(L_ACT1_8)*(0.075751)+V(L_ACT1_9)*(0.235079)+V(L_ACT1_10)*(0.080266)+V(L_ACT1_11)*(-0.034430)+V(L_ACT1_12)*(0.157573)+V(L_ACT1_13)*(0.133040)+V(L_ACT1_14)*(-0.018706)+V(L_ACT1_15)*(-0.119657)+V(L_ACT1_16)*(-0.097665)+V(L_ACT1_17)*(-0.171140)+V(L_ACT1_18)*(-0.066478)+V(L_ACT1_19)*(0.166309)+V(L_ACT1_20)*(0.124289)+V(L_ACT1_21)*(-0.146226)+V(L_ACT1_22)*(-0.162288)+V(L_ACT1_23)*(-0.214174)+V(L_ACT1_24)*(0.028281)+V(L_ACT1_25)*(-0.021645)+V(L_ACT1_26)*(-0.154146)+V(L_ACT1_27)*(-0.037620)+V(L_ACT1_28)*(-0.128024)+V(L_ACT1_29)*(-0.018993)+V(L_ACT1_30)*(-0.006736)+V(L_ACT1_31)*(0.002615)+V(L_ACT1_32)*(0.072705)+(0.088963))
B2_5 L2_5 0 V=(V(L_ACT1_1)*(-0.085566)+V(L_ACT1_2)*(-0.161670)+V(L_ACT1_3)*(-0.064274)+V(L_ACT1_4)*(-0.051710)+V(L_ACT1_5)*(0.001126)+V(L_ACT1_6)*(-0.152769)+V(L_ACT1_7)*(0.131411)+V(L_ACT1_8)*(-0.006619)+V(L_ACT1_9)*(0.098095)+V(L_ACT1_10)*(-0.107359)+V(L_ACT1_11)*(-0.068960)+V(L_ACT1_12)*(0.099391)+V(L_ACT1_13)*(-0.007186)+V(L_ACT1_14)*(0.036720)+V(L_ACT1_15)*(0.013167)+V(L_ACT1_16)*(0.098745)+V(L_ACT1_17)*(0.023342)+V(L_ACT1_18)*(-0.033140)+V(L_ACT1_19)*(0.093707)+V(L_ACT1_20)*(-0.166766)+V(L_ACT1_21)*(-0.088985)+V(L_ACT1_22)*(-0.107786)+V(L_ACT1_23)*(0.004567)+V(L_ACT1_24)*(-0.029251)+V(L_ACT1_25)*(-0.023790)+V(L_ACT1_26)*(0.210934)+V(L_ACT1_27)*(0.192894)+V(L_ACT1_28)*(-0.132524)+V(L_ACT1_29)*(0.096560)+V(L_ACT1_30)*(-0.066583)+V(L_ACT1_31)*(-0.163500)+V(L_ACT1_32)*(-0.000321)+(0.033796))
B2_6 L2_6 0 V=(V(L_ACT1_1)*(-0.088219)+V(L_ACT1_2)*(0.044367)+V(L_ACT1_3)*(-0.168456)+V(L_ACT1_4)*(0.148239)+V(L_ACT1_5)*(-0.206833)+V(L_ACT1_6)*(0.174220)+V(L_ACT1_7)*(0.015952)+V(L_ACT1_8)*(0.181608)+V(L_ACT1_9)*(0.185881)+V(L_ACT1_10)*(0.059591)+V(L_ACT1_11)*(0.027398)+V(L_ACT1_12)*(0.148863)+V(L_ACT1_13)*(-0.089213)+V(L_ACT1_14)*(0.168253)+V(L_ACT1_15)*(0.040729)+V(L_ACT1_16)*(-0.008860)+V(L_ACT1_17)*(0.000202)+V(L_ACT1_18)*(0.046574)+V(L_ACT1_19)*(-0.006837)+V(L_ACT1_20)*(0.077959)+V(L_ACT1_21)*(-0.036301)+V(L_ACT1_22)*(-0.005396)+V(L_ACT1_23)*(-0.147665)+V(L_ACT1_24)*(0.074566)+V(L_ACT1_25)*(-0.023581)+V(L_ACT1_26)*(0.090087)+V(L_ACT1_27)*(-0.122130)+V(L_ACT1_28)*(-0.209058)+V(L_ACT1_29)*(-0.066808)+V(L_ACT1_30)*(-0.201508)+V(L_ACT1_31)*(0.099076)+V(L_ACT1_32)*(-0.072489)+(0.214714))
B2_7 L2_7 0 V=(V(L_ACT1_1)*(-0.247854)+V(L_ACT1_2)*(0.004369)+V(L_ACT1_3)*(-0.135639)+V(L_ACT1_4)*(0.161874)+V(L_ACT1_5)*(-0.088220)+V(L_ACT1_6)*(0.006630)+V(L_ACT1_7)*(0.109624)+V(L_ACT1_8)*(0.118057)+V(L_ACT1_9)*(0.064634)+V(L_ACT1_10)*(0.022960)+V(L_ACT1_11)*(0.086487)+V(L_ACT1_12)*(-0.125074)+V(L_ACT1_13)*(-0.123218)+V(L_ACT1_14)*(0.119120)+V(L_ACT1_15)*(-0.042813)+V(L_ACT1_16)*(-0.058337)+V(L_ACT1_17)*(0.034485)+V(L_ACT1_18)*(0.188747)+V(L_ACT1_19)*(0.313836)+V(L_ACT1_20)*(-0.178550)+V(L_ACT1_21)*(-0.029320)+V(L_ACT1_22)*(0.037018)+V(L_ACT1_23)*(0.013945)+V(L_ACT1_24)*(0.130544)+V(L_ACT1_25)*(0.070187)+V(L_ACT1_26)*(-0.147673)+V(L_ACT1_27)*(0.054355)+V(L_ACT1_28)*(-0.098327)+V(L_ACT1_29)*(0.017908)+V(L_ACT1_30)*(-0.012014)+V(L_ACT1_31)*(0.076507)+V(L_ACT1_32)*(0.086757)+(0.168249))
B2_8 L2_8 0 V=(V(L_ACT1_1)*(-0.107527)+V(L_ACT1_2)*(0.163391)+V(L_ACT1_3)*(0.145092)+V(L_ACT1_4)*(-0.036676)+V(L_ACT1_5)*(-0.017167)+V(L_ACT1_6)*(-0.147841)+V(L_ACT1_7)*(-0.063868)+V(L_ACT1_8)*(-0.050353)+V(L_ACT1_9)*(0.056014)+V(L_ACT1_10)*(-0.056650)+V(L_ACT1_11)*(-0.059242)+V(L_ACT1_12)*(-0.151599)+V(L_ACT1_13)*(-0.065901)+V(L_ACT1_14)*(-0.173729)+V(L_ACT1_15)*(-0.158671)+V(L_ACT1_16)*(0.038431)+V(L_ACT1_17)*(-0.033088)+V(L_ACT1_18)*(0.108975)+V(L_ACT1_19)*(-0.120763)+V(L_ACT1_20)*(-0.094099)+V(L_ACT1_21)*(0.071462)+V(L_ACT1_22)*(0.155886)+V(L_ACT1_23)*(-0.049431)+V(L_ACT1_24)*(0.051098)+V(L_ACT1_25)*(0.032588)+V(L_ACT1_26)*(0.005487)+V(L_ACT1_27)*(-0.068877)+V(L_ACT1_28)*(0.107408)+V(L_ACT1_29)*(0.120071)+V(L_ACT1_30)*(-0.161360)+V(L_ACT1_31)*(0.012871)+V(L_ACT1_32)*(0.048241)+(-0.125543))
B2_9 L2_9 0 V=(V(L_ACT1_1)*(-0.207682)+V(L_ACT1_2)*(0.026251)+V(L_ACT1_3)*(-0.149401)+V(L_ACT1_4)*(0.172148)+V(L_ACT1_5)*(0.057006)+V(L_ACT1_6)*(0.185928)+V(L_ACT1_7)*(0.149295)+V(L_ACT1_8)*(-0.106970)+V(L_ACT1_9)*(0.240654)+V(L_ACT1_10)*(0.042982)+V(L_ACT1_11)*(0.020039)+V(L_ACT1_12)*(-0.049739)+V(L_ACT1_13)*(0.177462)+V(L_ACT1_14)*(0.033039)+V(L_ACT1_15)*(0.087235)+V(L_ACT1_16)*(-0.019519)+V(L_ACT1_17)*(0.133247)+V(L_ACT1_18)*(0.081042)+V(L_ACT1_19)*(0.141748)+V(L_ACT1_20)*(0.007413)+V(L_ACT1_21)*(0.090278)+V(L_ACT1_22)*(-0.001001)+V(L_ACT1_23)*(-0.132639)+V(L_ACT1_24)*(0.180537)+V(L_ACT1_25)*(-0.194263)+V(L_ACT1_26)*(-0.179916)+V(L_ACT1_27)*(-0.012737)+V(L_ACT1_28)*(-0.096658)+V(L_ACT1_29)*(0.176473)+V(L_ACT1_30)*(0.125035)+V(L_ACT1_31)*(0.183419)+V(L_ACT1_32)*(-0.131586)+(-0.055426))
B2_10 L2_10 0 V=(V(L_ACT1_1)*(0.223489)+V(L_ACT1_2)*(-0.000175)+V(L_ACT1_3)*(0.014489)+V(L_ACT1_4)*(-0.116280)+V(L_ACT1_5)*(-0.052792)+V(L_ACT1_6)*(0.061171)+V(L_ACT1_7)*(-0.011171)+V(L_ACT1_8)*(-0.139987)+V(L_ACT1_9)*(-0.036964)+V(L_ACT1_10)*(-0.006463)+V(L_ACT1_11)*(-0.044069)+V(L_ACT1_12)*(0.173242)+V(L_ACT1_13)*(-0.100474)+V(L_ACT1_14)*(-0.078123)+V(L_ACT1_15)*(0.063941)+V(L_ACT1_16)*(0.066554)+V(L_ACT1_17)*(-0.165293)+V(L_ACT1_18)*(-0.190369)+V(L_ACT1_19)*(-0.192562)+V(L_ACT1_20)*(-0.026011)+V(L_ACT1_21)*(-0.021673)+V(L_ACT1_22)*(0.065118)+V(L_ACT1_23)*(-0.013335)+V(L_ACT1_24)*(0.013964)+V(L_ACT1_25)*(0.116939)+V(L_ACT1_26)*(-0.033918)+V(L_ACT1_27)*(0.240118)+V(L_ACT1_28)*(0.383603)+V(L_ACT1_29)*(0.047262)+V(L_ACT1_30)*(-0.055522)+V(L_ACT1_31)*(-0.113439)+V(L_ACT1_32)*(0.058572)+(0.083639))
B2_11 L2_11 0 V=(V(L_ACT1_1)*(-0.054570)+V(L_ACT1_2)*(0.206599)+V(L_ACT1_3)*(-0.189172)+V(L_ACT1_4)*(0.153111)+V(L_ACT1_5)*(-0.119552)+V(L_ACT1_6)*(0.115081)+V(L_ACT1_7)*(0.007588)+V(L_ACT1_8)*(-0.045404)+V(L_ACT1_9)*(0.141949)+V(L_ACT1_10)*(0.090675)+V(L_ACT1_11)*(-0.188620)+V(L_ACT1_12)*(0.012502)+V(L_ACT1_13)*(-0.044611)+V(L_ACT1_14)*(0.124062)+V(L_ACT1_15)*(-0.096107)+V(L_ACT1_16)*(-0.019447)+V(L_ACT1_17)*(0.080325)+V(L_ACT1_18)*(-0.045095)+V(L_ACT1_19)*(0.084980)+V(L_ACT1_20)*(0.060885)+V(L_ACT1_21)*(-0.095061)+V(L_ACT1_22)*(-0.093897)+V(L_ACT1_23)*(0.015229)+V(L_ACT1_24)*(0.113783)+V(L_ACT1_25)*(0.059669)+V(L_ACT1_26)*(0.047108)+V(L_ACT1_27)*(0.009032)+V(L_ACT1_28)*(-0.130136)+V(L_ACT1_29)*(0.107264)+V(L_ACT1_30)*(0.026690)+V(L_ACT1_31)*(-0.134274)+V(L_ACT1_32)*(-0.107955)+(0.183581))
B2_12 L2_12 0 V=(V(L_ACT1_1)*(-0.164015)+V(L_ACT1_2)*(0.147398)+V(L_ACT1_3)*(-0.187345)+V(L_ACT1_4)*(0.017702)+V(L_ACT1_5)*(-0.100462)+V(L_ACT1_6)*(0.107591)+V(L_ACT1_7)*(0.145380)+V(L_ACT1_8)*(0.003259)+V(L_ACT1_9)*(0.207910)+V(L_ACT1_10)*(0.072773)+V(L_ACT1_11)*(0.009481)+V(L_ACT1_12)*(0.148508)+V(L_ACT1_13)*(-0.032846)+V(L_ACT1_14)*(-0.007049)+V(L_ACT1_15)*(-0.111063)+V(L_ACT1_16)*(-0.023724)+V(L_ACT1_17)*(-0.083978)+V(L_ACT1_18)*(0.003028)+V(L_ACT1_19)*(0.171713)+V(L_ACT1_20)*(-0.123234)+V(L_ACT1_21)*(0.067038)+V(L_ACT1_22)*(-0.073486)+V(L_ACT1_23)*(-0.073370)+V(L_ACT1_24)*(-0.036068)+V(L_ACT1_25)*(0.107316)+V(L_ACT1_26)*(0.144961)+V(L_ACT1_27)*(0.067312)+V(L_ACT1_28)*(-0.155623)+V(L_ACT1_29)*(0.135569)+V(L_ACT1_30)*(0.134752)+V(L_ACT1_31)*(0.141936)+V(L_ACT1_32)*(0.072811)+(-0.116490))
B2_13 L2_13 0 V=(V(L_ACT1_1)*(0.114476)+V(L_ACT1_2)*(-0.027405)+V(L_ACT1_3)*(-0.052727)+V(L_ACT1_4)*(0.065683)+V(L_ACT1_5)*(0.166178)+V(L_ACT1_6)*(-0.142116)+V(L_ACT1_7)*(0.091474)+V(L_ACT1_8)*(0.072936)+V(L_ACT1_9)*(-0.161924)+V(L_ACT1_10)*(0.140854)+V(L_ACT1_11)*(0.136692)+V(L_ACT1_12)*(0.127709)+V(L_ACT1_13)*(0.144877)+V(L_ACT1_14)*(-0.026892)+V(L_ACT1_15)*(0.131950)+V(L_ACT1_16)*(0.115149)+V(L_ACT1_17)*(0.108755)+V(L_ACT1_18)*(0.032665)+V(L_ACT1_19)*(-0.182522)+V(L_ACT1_20)*(0.185729)+V(L_ACT1_21)*(-0.099219)+V(L_ACT1_22)*(-0.113606)+V(L_ACT1_23)*(0.143149)+V(L_ACT1_24)*(-0.096476)+V(L_ACT1_25)*(0.207408)+V(L_ACT1_26)*(-0.077965)+V(L_ACT1_27)*(0.167008)+V(L_ACT1_28)*(0.377073)+V(L_ACT1_29)*(-0.097539)+V(L_ACT1_30)*(-0.000180)+V(L_ACT1_31)*(-0.093315)+V(L_ACT1_32)*(0.066650)+(0.057935))
B2_14 L2_14 0 V=(V(L_ACT1_1)*(0.018004)+V(L_ACT1_2)*(0.107695)+V(L_ACT1_3)*(-0.049562)+V(L_ACT1_4)*(0.056062)+V(L_ACT1_5)*(-0.148161)+V(L_ACT1_6)*(-0.055862)+V(L_ACT1_7)*(-0.033320)+V(L_ACT1_8)*(-0.097387)+V(L_ACT1_9)*(-0.101050)+V(L_ACT1_10)*(0.063677)+V(L_ACT1_11)*(0.070553)+V(L_ACT1_12)*(0.003701)+V(L_ACT1_13)*(-0.150393)+V(L_ACT1_14)*(0.098320)+V(L_ACT1_15)*(0.156894)+V(L_ACT1_16)*(0.167964)+V(L_ACT1_17)*(-0.059994)+V(L_ACT1_18)*(-0.163817)+V(L_ACT1_19)*(0.052296)+V(L_ACT1_20)*(-0.005426)+V(L_ACT1_21)*(0.035216)+V(L_ACT1_22)*(-0.017463)+V(L_ACT1_23)*(-0.016595)+V(L_ACT1_24)*(-0.204541)+V(L_ACT1_25)*(-0.092124)+V(L_ACT1_26)*(-0.009211)+V(L_ACT1_27)*(0.130601)+V(L_ACT1_28)*(-0.039495)+V(L_ACT1_29)*(-0.143474)+V(L_ACT1_30)*(0.217161)+V(L_ACT1_31)*(-0.078605)+V(L_ACT1_32)*(0.002884)+(-0.091448))
B2_15 L2_15 0 V=(V(L_ACT1_1)*(-0.036585)+V(L_ACT1_2)*(0.063880)+V(L_ACT1_3)*(-0.095808)+V(L_ACT1_4)*(0.152895)+V(L_ACT1_5)*(-0.158315)+V(L_ACT1_6)*(0.060939)+V(L_ACT1_7)*(0.155177)+V(L_ACT1_8)*(0.081892)+V(L_ACT1_9)*(-0.012924)+V(L_ACT1_10)*(0.121594)+V(L_ACT1_11)*(-0.111990)+V(L_ACT1_12)*(0.068933)+V(L_ACT1_13)*(0.037151)+V(L_ACT1_14)*(-0.088725)+V(L_ACT1_15)*(0.121770)+V(L_ACT1_16)*(0.110838)+V(L_ACT1_17)*(0.025722)+V(L_ACT1_18)*(0.005027)+V(L_ACT1_19)*(0.162684)+V(L_ACT1_20)*(-0.128752)+V(L_ACT1_21)*(0.058296)+V(L_ACT1_22)*(0.082818)+V(L_ACT1_23)*(-0.186276)+V(L_ACT1_24)*(-0.023189)+V(L_ACT1_25)*(-0.042188)+V(L_ACT1_26)*(-0.105368)+V(L_ACT1_27)*(-0.016288)+V(L_ACT1_28)*(-0.364140)+V(L_ACT1_29)*(-0.054458)+V(L_ACT1_30)*(0.120978)+V(L_ACT1_31)*(0.098662)+V(L_ACT1_32)*(-0.070980)+(-0.063668))
B2_16 L2_16 0 V=(V(L_ACT1_1)*(0.094816)+V(L_ACT1_2)*(-0.045166)+V(L_ACT1_3)*(-0.131735)+V(L_ACT1_4)*(-0.035818)+V(L_ACT1_5)*(0.071727)+V(L_ACT1_6)*(-0.025802)+V(L_ACT1_7)*(-0.157183)+V(L_ACT1_8)*(-0.091544)+V(L_ACT1_9)*(0.083832)+V(L_ACT1_10)*(-0.026725)+V(L_ACT1_11)*(-0.111142)+V(L_ACT1_12)*(-0.093134)+V(L_ACT1_13)*(0.074923)+V(L_ACT1_14)*(-0.069976)+V(L_ACT1_15)*(-0.012169)+V(L_ACT1_16)*(-0.022156)+V(L_ACT1_17)*(-0.143369)+V(L_ACT1_18)*(-0.019001)+V(L_ACT1_19)*(0.170430)+V(L_ACT1_20)*(-0.007040)+V(L_ACT1_21)*(-0.052095)+V(L_ACT1_22)*(0.012571)+V(L_ACT1_23)*(-0.001956)+V(L_ACT1_24)*(-0.070479)+V(L_ACT1_25)*(0.188493)+V(L_ACT1_26)*(0.111832)+V(L_ACT1_27)*(-0.078504)+V(L_ACT1_28)*(-0.024308)+V(L_ACT1_29)*(-0.072603)+V(L_ACT1_30)*(-0.083016)+V(L_ACT1_31)*(0.133637)+V(L_ACT1_32)*(-0.004464)+(0.032121))
* ACTIVATION LAYER 2: RELU
B_ACT2_1 L_ACT2_1 0 V=(IF(V(L2_1)>0,V(L2_1),0))
B_ACT2_2 L_ACT2_2 0 V=(IF(V(L2_2)>0,V(L2_2),0))
B_ACT2_3 L_ACT2_3 0 V=(IF(V(L2_3)>0,V(L2_3),0))
B_ACT2_4 L_ACT2_4 0 V=(IF(V(L2_4)>0,V(L2_4),0))
B_ACT2_5 L_ACT2_5 0 V=(IF(V(L2_5)>0,V(L2_5),0))
B_ACT2_6 L_ACT2_6 0 V=(IF(V(L2_6)>0,V(L2_6),0))
B_ACT2_7 L_ACT2_7 0 V=(IF(V(L2_7)>0,V(L2_7),0))
B_ACT2_8 L_ACT2_8 0 V=(IF(V(L2_8)>0,V(L2_8),0))
B_ACT2_9 L_ACT2_9 0 V=(IF(V(L2_9)>0,V(L2_9),0))
B_ACT2_10 L_ACT2_10 0 V=(IF(V(L2_10)>0,V(L2_10),0))
B_ACT2_11 L_ACT2_11 0 V=(IF(V(L2_11)>0,V(L2_11),0))
B_ACT2_12 L_ACT2_12 0 V=(IF(V(L2_12)>0,V(L2_12),0))
B_ACT2_13 L_ACT2_13 0 V=(IF(V(L2_13)>0,V(L2_13),0))
B_ACT2_14 L_ACT2_14 0 V=(IF(V(L2_14)>0,V(L2_14),0))
B_ACT2_15 L_ACT2_15 0 V=(IF(V(L2_15)>0,V(L2_15),0))
B_ACT2_16 L_ACT2_16 0 V=(IF(V(L2_16)>0,V(L2_16),0))
* LAYER 3: LINEAR
B3_1 L3_1 0 V=(V(L_ACT2_1)*(0.105320)+V(L_ACT2_2)*(-0.356847)+V(L_ACT2_3)*(-0.290122)+V(L_ACT2_4)*(0.099256)+V(L_ACT2_5)*(-0.190800)+V(L_ACT2_6)*(0.245422)+V(L_ACT2_7)*(0.181454)+V(L_ACT2_8)*(-0.020837)+V(L_ACT2_9)*(0.234329)+V(L_ACT2_10)*(-0.365517)+V(L_ACT2_11)*(0.209686)+V(L_ACT2_12)*(0.242298)+V(L_ACT2_13)*(-0.130089)+V(L_ACT2_14)*(-0.272604)+V(L_ACT2_15)*(0.354239)+V(L_ACT2_16)*(-0.232107)+(-0.140361))
* ACTIVATION LAYER 3: RELU
B_ACT3_1 L_ACT3_1 0 V=(IF(V(L3_1)>0,V(L3_1),0))
* Connect final internal node L_ACT3_1 to external output NNOUT1
B_OUT NNOUT1 0 V=V(L_ACT3_1)
.ENDS ActorSubckt